`timescale 1ns / 1ps
module adder( input [31:0] inp , output wire [31:0] out
    );

        assign out = inp + 1  ;

endmodule
