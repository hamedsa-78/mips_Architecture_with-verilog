`timescale 1ns / 1ps
module ALU_control(
input [1:0]ALU_op,
input [5:0]inst,
output reg [3:0]op,
output reg JR
 );
 
always @(*)
begin
JR = 0 ; 
	if(ALU_op == 2'b00)
	begin
	op = 4'b0010 ;
	end
	else if(ALU_op == 2'b01)
	begin
	op = 4'b0110 ;
	end
	else if(ALU_op == 2'b10)
	begin
		if(inst == 6'b100000)
		begin
		op = 4'b0010 ;
		end
		if(inst == 6'b011000)
		begin
		op = 4'b0010 ;
		end
		if(inst == 6'b100010)
		begin
		op = 4'b0110 ;
		end
		if(inst == 6'b100100)
		begin 
		op = 4'b0000 ;
		end
		if(inst == 6'b100101)
		begin
		op = 4'b0001 ;
		end
		if(inst == 6'b101010)
		begin
		op = 4'b0111 ;
		end
		if(inst == 6'b001100)//andi
		begin
		op = 4'b0000 ;
		end
		if(inst == 6'b001101)//ori
		begin
		op = 4'b0001 ;
		end
		
		if(inst == 6'b001000)//JR
		begin
		JR = 1 ;
		op = 4'b0011 ;
		end
		
	end
end


endmodule
